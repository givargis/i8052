-- sqrt.hex
-- Wed Jul 16 07:58:05 2025

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_ARITH.all;

use WORK.I8052_PKG.all;

entity I8052_ROM is
  port(rst : in  STD_LOGIC;
       clk : in  STD_LOGIC;
       addr: in  UNSIGNED (11 downto 0);
       data: out UNSIGNED (7 downto 0);
       rd  : in  STD_LOGIC);
end I8052_ROM;

architecture BEHAVIORAL of I8052_ROM is
  type ROM_TYPE is array (0 to 2132) of UNSIGNED (7 downto 0);
  constant PROGRAM : ROM_TYPE := (
    "00000010",  -- 00000: LJMP
    "00000000",
    "01001100",
    "00000000",  -- 00003: NOP
    "00000000",  -- 00004: NOP
    "00000000",  -- 00005: NOP
    "00000000",  -- 00006: NOP
    "00000000",  -- 00007: NOP
    "00000000",  -- 00008: NOP
    "00000000",  -- 00009: NOP
    "11100010",  -- 00010: MOVX_1
    "11111011",  -- 00011: MOV_5
    "11101010",  -- 00012: MOV_1
    "11110010",  -- 00013: MOVX_3
    "10000000",  -- 00014: SJMP
    "00101100",
    "00000000",  -- 00016: NOP
    "00000000",  -- 00017: NOP
    "11100000",  -- 00018: MOVX_2
    "11111011",  -- 00019: MOV_5
    "11101010",  -- 00020: MOV_1
    "11110000",  -- 00021: MOVX_4
    "10000000",  -- 00022: SJMP
    "00100100",
    "11100110",  -- 00024: MOV_3
    "10110101",  -- 00025: CJNE_1
    "00000010",
    "00000010",
    "11101011",  -- 00028: MOV_1
    "11110110",  -- 00029: MOV_13
    "00100010",  -- 00030: RET
    "00000000",  -- 00031: NOP
    "11100010",  -- 00032: MOVX_1
    "10110101",  -- 00033: CJNE_1
    "00000010",
    "00000010",
    "11101011",  -- 00036: MOV_1
    "11110010",  -- 00037: MOVX_3
    "00100010",  -- 00038: RET
    "00000000",  -- 00039: NOP
    "11100000",  -- 00040: MOVX_2
    "10110101",  -- 00041: CJNE_1
    "00000010",
    "00000010",
    "11101011",  -- 00044: MOV_1
    "11110000",  -- 00045: MOVX_4
    "00100010",  -- 00046: RET
    "00110000",  -- 00047: JNB
    "11110110",
    "11100000",
    "10101000",  -- 00050: MOV_6
    "10000010",
    "00100000",  -- 00052: JB
    "11110101",
    "11010011",
    "11101010",  -- 00055: MOV_1
    "11000110",  -- 00056: XCH_3
    "11110101",  -- 00057: MOV_8
    "10000010",
    "00100010",  -- 00059: RET
    "10001011",  -- 00060: MOV_9
    "10000010",
    "00100010",  -- 00062: RET
    "00110000",  -- 00063: JNB
    "11110110",
    "11100110",
    "10101000",  -- 00066: MOV_6
    "10000010",
    "00100000",  -- 00068: JB
    "11110101",
    "11011001",
    "10000000",  -- 00071: SJMP
    "11001111",
    "00000010",  -- 00073: LJMP
    "00000000",
    "10101000",
    "01110101",  -- 00076: MOV_12
    "10000001",
    "00010101",
    "00010010",  -- 00079: LCALL
    "00001000",
    "00111101",
    "11100101",  -- 00082: MOV_2
    "10000010",
    "01100000",  -- 00084: JZ
    "00000011",
    "00000010",  -- 00086: LJMP
    "00000000",
    "01001001",
    "01111001",  -- 00089: MOV_7
    "00000000",
    "11101001",  -- 00091: MOV_1
    "01000100",  -- 00092: ORL_4
    "00000000",
    "01100000",  -- 00094: JZ
    "00011011",
    "01111010",  -- 00096: MOV_7
    "00000000",
    "10010000",  -- 00098: MOV_18
    "00001000",
    "01010011",
    "01111000",  -- 00101: MOV_7
    "00000001",
    "01110101",  -- 00103: MOV_12
    "10100000",
    "00000000",
    "11100100",  -- 00106: CLR_1
    "10010011",  -- 00107: MOVC_1
    "11110010",  -- 00108: MOVX_3
    "10100011",  -- 00109: INC_5
    "00001000",  -- 00110: INC_2
    "10111000",  -- 00111: CJNE_3
    "00000000",
    "00000010",
    "00000101",  -- 00114: INC_3
    "10100000",
    "11011001",  -- 00116: DJNZ_1
    "11110100",
    "11011010",  -- 00118: DJNZ_1
    "11110010",
    "01110101",  -- 00120: MOV_12
    "10100000",
    "11111111",
    "11100100",  -- 00123: CLR_1
    "01111000",  -- 00124: MOV_7
    "11111111",
    "11110110",  -- 00126: MOV_13
    "11011000",  -- 00127: DJNZ_1
    "11111101",
    "01111000",  -- 00129: MOV_7
    "00000000",
    "11101000",  -- 00131: MOV_1
    "01000100",  -- 00132: ORL_4
    "00000000",
    "01100000",  -- 00134: JZ
    "00001010",
    "01111001",  -- 00136: MOV_7
    "00000001",
    "01110101",  -- 00138: MOV_12
    "10100000",
    "00000000",
    "11100100",  -- 00141: CLR_1
    "11110011",  -- 00142: MOVX_3
    "00001001",  -- 00143: INC_2
    "11011000",  -- 00144: DJNZ_1
    "11111100",
    "01111000",  -- 00146: MOV_7
    "00000000",
    "11101000",  -- 00148: MOV_1
    "01000100",  -- 00149: ORL_4
    "00000000",
    "01100000",  -- 00151: JZ
    "00001100",
    "01111001",  -- 00153: MOV_7
    "00000000",
    "10010000",  -- 00155: MOV_18
    "00000000",
    "00000001",
    "11100100",  -- 00158: CLR_1
    "11110000",  -- 00159: MOVX_4
    "10100011",  -- 00160: INC_5
    "11011000",  -- 00161: DJNZ_1
    "11111100",
    "11011001",  -- 00163: DJNZ_1
    "11111010",
    "00000010",  -- 00165: LJMP
    "00000000",
    "01001001",
    "01110101",  -- 00168: MOV_12
    "10000000",
    "00001001",
    "01110101",  -- 00171: MOV_12
    "10010000",
    "00010000",
    "01110101",  -- 00174: MOV_12
    "10100000",
    "00011001",
    "10010000",  -- 00177: MOV_18
    "00000000",
    "00000000",
    "01110101",  -- 00180: MOV_12
    "11110000",
    "11001000",
    "01110100",  -- 00183: MOV_4
    "01000001",
    "00010010",  -- 00185: LCALL
    "00000000",
    "11000100",
    "00010010",  -- 00188: LCALL
    "00000110",
    "01100011",
    "10000101",  -- 00191: MOV_10
    "10000010",
    "10110000",
    "10000000",  -- 00194: SJMP
    "11111110",
    "11000000",  -- 00196: PUSH
    "00001000",
    "10000101",  -- 00198: MOV_10
    "10000001",
    "00001000",
    "10101100",  -- 00201: MOV_6
    "10000010",
    "10101101",  -- 00203: MOV_6
    "10000011",
    "10101110",  -- 00205: MOV_6
    "11110000",
    "11111111",  -- 00207: MOV_5
    "11100101",  -- 00208: MOV_2
    "10000001",
    "00100100",  -- 00210: ADD_4
    "00001010",
    "11110101",  -- 00212: MOV_8
    "10000001",
    "10001100",  -- 00214: MOV_9
    "11110000",
    "11101101",  -- 00216: MOV_1
    "01000010",  -- 00217: ORL_5
    "11110000",
    "11101110",  -- 00219: MOV_1
    "01000010",  -- 00220: ORL_5
    "11110000",
    "11101111",  -- 00222: MOV_1
    "01010100",  -- 00223: ANL_4
    "01111111",
    "01000101",  -- 00225: ORL_2
    "11110000",
    "01110000",  -- 00227: JNZ
    "00001010",
    "10001100",  -- 00229: MOV_9
    "10000010",
    "10001101",  -- 00231: MOV_9
    "10000011",
    "10001110",  -- 00233: MOV_9
    "11110000",
    "11101111",  -- 00235: MOV_1
    "00000010",  -- 00236: LJMP
    "00000011",
    "00001101",
    "11000000",  -- 00239: PUSH
    "00000111",
    "11000000",  -- 00241: PUSH
    "00000110",
    "11000000",  -- 00243: PUSH
    "00000101",
    "11000000",  -- 00245: PUSH
    "00000100",
    "11100100",  -- 00247: CLR_1
    "11000000",  -- 00248: PUSH
    "11100000",
    "11000000",  -- 00250: PUSH
    "11100000",
    "01110100",  -- 00252: MOV_4
    "10000000",
    "11000000",  -- 00254: PUSH
    "11100000",
    "01110100",  -- 00256: MOV_4
    "00111111",
    "11000000",  -- 00258: PUSH
    "11100000",
    "10001100",  -- 00260: MOV_9
    "10000010",
    "10001101",  -- 00262: MOV_9
    "10000011",
    "10001110",  -- 00264: MOV_9
    "11110000",
    "11101111",  -- 00266: MOV_1
    "00010010",  -- 00267: LCALL
    "00000111",
    "11101010",
    "10101011",  -- 00270: MOV_6
    "10000010",
    "11100101",  -- 00272: MOV_2
    "10000001",
    "00100100",  -- 00274: ADD_4
    "11111100",
    "11110101",  -- 00276: MOV_8
    "10000001",
    "11010000",  -- 00278: POP
    "00000100",
    "11010000",  -- 00280: POP
    "00000101",
    "11010000",  -- 00282: POP
    "00000110",
    "11010000",  -- 00284: POP
    "00000111",
    "11101011",  -- 00286: MOV_1
    "01100000",  -- 00287: JZ
    "00001011",
    "10010000",  -- 00289: MOV_18
    "00000000",
    "00000000",
    "01110101",  -- 00292: MOV_12
    "11110000",
    "10000000",
    "01110100",  -- 00295: MOV_4
    "00111111",
    "00000010",  -- 00297: LJMP
    "00000011",
    "00001101",
    "11000000",  -- 00300: PUSH
    "00000111",
    "11000000",  -- 00302: PUSH
    "00000110",
    "11000000",  -- 00304: PUSH
    "00000101",
    "11000000",  -- 00306: PUSH
    "00000100",
    "11100100",  -- 00308: CLR_1
    "11000000",  -- 00309: PUSH
    "11100000",
    "11000000",  -- 00311: PUSH
    "11100000",
    "11000000",  -- 00313: PUSH
    "11100000",
    "11000000",  -- 00315: PUSH
    "11100000",
    "10001100",  -- 00317: MOV_9
    "10000010",
    "10001101",  -- 00319: MOV_9
    "10000011",
    "10001110",  -- 00321: MOV_9
    "11110000",
    "11101111",  -- 00323: MOV_1
    "00010010",  -- 00324: LCALL
    "00000011",
    "00010011",
    "10101011",  -- 00327: MOV_6
    "10000010",
    "11100101",  -- 00329: MOV_2
    "10000001",
    "00100100",  -- 00331: ADD_4
    "11111100",
    "11110101",  -- 00333: MOV_8
    "10000001",
    "11010000",  -- 00335: POP
    "00000100",
    "11010000",  -- 00337: POP
    "00000101",
    "11010000",  -- 00339: POP
    "00000110",
    "11010000",  -- 00341: POP
    "00000111",
    "11101011",  -- 00343: MOV_1
    "01100000",  -- 00344: JZ
    "00001111",
    "01110101",  -- 00346: MOV_12
    "00001001",
    "00100001",
    "01110101",  -- 00349: MOV_12
    "00001010",
    "00000000",
    "10010000",  -- 00352: MOV_18
    "00000000",
    "00000000",
    "11100100",  -- 00355: CLR_1
    "11110101",  -- 00356: MOV_8
    "11110000",
    "00000010",  -- 00358: LJMP
    "00000011",
    "00001101",
    "11100101",  -- 00361: MOV_2
    "00001000",
    "00100100",  -- 00363: ADD_4
    "00001001",
    "11110101",  -- 00365: MOV_8
    "00001011",
    "01110101",  -- 00367: MOV_12
    "00001100",
    "00000000",
    "01110101",  -- 00370: MOV_12
    "00001101",
    "01000000",
    "10001100",  -- 00373: MOV_9
    "10000010",
    "10001101",  -- 00375: MOV_9
    "10000011",
    "10001110",  -- 00377: MOV_9
    "11110000",
    "11101111",  -- 00379: MOV_1
    "00010010",  -- 00380: LCALL
    "00000100",
    "10100010",
    "11001000",  -- 00383: XCH_1
    "11100101",  -- 00384: MOV_2
    "00001000",
    "00100100",  -- 00386: ADD_4
    "00000101",
    "11001000",  -- 00388: XCH_1
    "10100110",  -- 00389: MOV_14
    "10000010",
    "00001000",  -- 00391: INC_2
    "10100110",  -- 00392: MOV_14
    "10000011",
    "00001000",  -- 00394: INC_2
    "10100110",  -- 00395: MOV_14
    "11110000",
    "00001000",  -- 00397: INC_2
    "11110110",  -- 00398: MOV_13
    "11100101",  -- 00399: MOV_2
    "00001000",
    "00100100",  -- 00401: ADD_4
    "00000101",
    "11111000",  -- 00403: MOV_5
    "11100110",  -- 00404: MOV_3
    "11000000",  -- 00405: PUSH
    "11100000",
    "00001000",  -- 00407: INC_2
    "11100110",  -- 00408: MOV_3
    "11000000",  -- 00409: PUSH
    "11100000",
    "00001000",  -- 00411: INC_2
    "11100110",  -- 00412: MOV_3
    "11000000",  -- 00413: PUSH
    "11100000",
    "00001000",  -- 00415: INC_2
    "11100110",  -- 00416: MOV_3
    "11000000",  -- 00417: PUSH
    "11100000",
    "10010000",  -- 00419: MOV_18
    "00010100",
    "10111010",
    "01110101",  -- 00422: MOV_12
    "11110000",
    "00010111",
    "01110100",  -- 00425: MOV_4
    "00111111",
    "00010010",  -- 00427: LCALL
    "00000110",
    "10100011",
    "10101010",  -- 00430: MOV_6
    "10000010",
    "10101011",  -- 00432: MOV_6
    "10000011",
    "10101110",  -- 00434: MOV_6
    "11110000",
    "11111111",  -- 00436: MOV_5
    "11100101",  -- 00437: MOV_2
    "10000001",
    "00100100",  -- 00439: ADD_4
    "11111100",
    "11110101",  -- 00441: MOV_8
    "10000001",
    "01110100",  -- 00443: MOV_4
    "10101000",
    "11000000",  -- 00445: PUSH
    "11100000",
    "00000100",  -- 00447: INC_1
    "11000000",  -- 00448: PUSH
    "11100000",
    "01110100",  -- 00450: MOV_4
    "11010101",
    "11000000",  -- 00452: PUSH
    "11100000",
    "01110100",  -- 00454: MOV_4
    "00111110",
    "11000000",  -- 00456: PUSH
    "11100000",
    "10001010",  -- 00458: MOV_9
    "10000010",
    "10001011",  -- 00460: MOV_9
    "10000011",
    "10001110",  -- 00462: MOV_9
    "11110000",
    "11101111",  -- 00464: MOV_1
    "00010010",  -- 00465: LCALL
    "00000011",
    "01000011",
    "10101000",  -- 00468: MOV_6
    "00001000",
    "00001000",  -- 00470: INC_2
    "10100110",  -- 00471: MOV_14
    "10000010",
    "00001000",  -- 00473: INC_2
    "10100110",  -- 00474: MOV_14
    "10000011",
    "00001000",  -- 00476: INC_2
    "10100110",  -- 00477: MOV_14
    "11110000",
    "00001000",  -- 00479: INC_2
    "11110110",  -- 00480: MOV_13
    "11100101",  -- 00481: MOV_2
    "10000001",
    "00100100",  -- 00483: ADD_4
    "11111100",
    "11110101",  -- 00485: MOV_8
    "10000001",
    "10101000",  -- 00487: MOV_6
    "00001000",
    "00001000",  -- 00489: INC_2
    "11100110",  -- 00490: MOV_3
    "11000000",  -- 00491: PUSH
    "11100000",
    "00001000",  -- 00493: INC_2
    "11100110",  -- 00494: MOV_3
    "11000000",  -- 00495: PUSH
    "11100000",
    "00001000",  -- 00497: INC_2
    "11100110",  -- 00498: MOV_3
    "11000000",  -- 00499: PUSH
    "11100000",
    "00001000",  -- 00501: INC_2
    "11100110",  -- 00502: MOV_3
    "11000000",  -- 00503: PUSH
    "11100000",
    "11100101",  -- 00505: MOV_2
    "00001000",
    "00100100",  -- 00507: ADD_4
    "00000101",
    "11111000",  -- 00509: MOV_5
    "10000110",  -- 00510: MOV_11
    "10000010",
    "00001000",  -- 00512: INC_2
    "10000110",  -- 00513: MOV_11
    "10000011",
    "00001000",  -- 00515: INC_2
    "10000110",  -- 00516: MOV_11
    "11110000",
    "00001000",  -- 00518: INC_2
    "11100110",  -- 00519: MOV_3
    "00010010",  -- 00520: LCALL
    "00000101",
    "10100000",
    "10101010",  -- 00523: MOV_6
    "10000010",
    "10101011",  -- 00525: MOV_6
    "10000011",
    "10101110",  -- 00527: MOV_6
    "11110000",
    "11111111",  -- 00529: MOV_5
    "11100101",  -- 00530: MOV_2
    "10000001",
    "00100100",  -- 00532: ADD_4
    "11111100",
    "11110101",  -- 00534: MOV_8
    "10000001",
    "11000000",  -- 00536: PUSH
    "00000010",
    "11000000",  -- 00538: PUSH
    "00000011",
    "11000000",  -- 00540: PUSH
    "00000110",
    "11000000",  -- 00542: PUSH
    "00000111",
    "10101000",  -- 00544: MOV_6
    "00001000",
    "00001000",  -- 00546: INC_2
    "10000110",  -- 00547: MOV_11
    "10000010",
    "00001000",  -- 00549: INC_2
    "10000110",  -- 00550: MOV_11
    "10000011",
    "00001000",  -- 00552: INC_2
    "10000110",  -- 00553: MOV_11
    "11110000",
    "00001000",  -- 00555: INC_2
    "11100110",  -- 00556: MOV_3
    "00010010",  -- 00557: LCALL
    "00000011",
    "01000011",
    "10101111",  -- 00560: MOV_6
    "10000010",
    "10101110",  -- 00562: MOV_6
    "10000011",
    "10101101",  -- 00564: MOV_6
    "11110000",
    "11111100",  -- 00566: MOV_5
    "11100101",  -- 00567: MOV_2
    "10000001",
    "00100100",  -- 00569: ADD_4
    "11111100",
    "11110101",  -- 00571: MOV_8
    "10000001",
    "01110101",  -- 00573: MOV_12
    "00001011",
    "11111110",
    "01110101",  -- 00576: MOV_12
    "00001100",
    "11111111",
    "10001111",  -- 00579: MOV_9
    "10000010",
    "10001110",  -- 00581: MOV_9
    "10000011",
    "10001101",  -- 00583: MOV_9
    "11110000",
    "11101100",  -- 00585: MOV_1
    "11000000",  -- 00586: PUSH
    "00000111",
    "11000000",  -- 00588: PUSH
    "00000110",
    "11000000",  -- 00590: PUSH
    "00000101",
    "11000000",  -- 00592: PUSH
    "00000100",
    "00010010",  -- 00594: LCALL
    "00000011",
    "11000101",
    "10101000",  -- 00597: MOV_6
    "00001000",
    "00001000",  -- 00599: INC_2
    "10100110",  -- 00600: MOV_14
    "10000010",
    "00001000",  -- 00602: INC_2
    "10100110",  -- 00603: MOV_14
    "10000011",
    "00001000",  -- 00605: INC_2
    "10100110",  -- 00606: MOV_14
    "11110000",
    "00001000",  -- 00608: INC_2
    "11110110",  -- 00609: MOV_13
    "11100101",  -- 00610: MOV_2
    "00001000",
    "00100100",  -- 00612: ADD_4
    "00000101",
    "11111000",  -- 00614: MOV_5
    "10000110",  -- 00615: MOV_11
    "10000010",
    "00001000",  -- 00617: INC_2
    "10000110",  -- 00618: MOV_11
    "10000011",
    "00001000",  -- 00620: INC_2
    "10000110",  -- 00621: MOV_11
    "11110000",
    "00001000",  -- 00623: INC_2
    "11100110",  -- 00624: MOV_3
    "00010010",  -- 00625: LCALL
    "00000101",
    "10100000",
    "10101100",  -- 00628: MOV_6
    "10000010",
    "10101101",  -- 00630: MOV_6
    "10000011",
    "10101110",  -- 00632: MOV_6
    "11110000",
    "11111111",  -- 00634: MOV_5
    "11100101",  -- 00635: MOV_2
    "10000001",
    "00100100",  -- 00637: ADD_4
    "11111100",
    "11110101",  -- 00639: MOV_8
    "10000001",
    "11000000",  -- 00641: PUSH
    "00000100",
    "11000000",  -- 00643: PUSH
    "00000101",
    "11000000",  -- 00645: PUSH
    "00000110",
    "11000000",  -- 00647: PUSH
    "00000111",
    "10101000",  -- 00649: MOV_6
    "00001000",
    "00001000",  -- 00651: INC_2
    "10000110",  -- 00652: MOV_11
    "10000010",
    "00001000",  -- 00654: INC_2
    "10000110",  -- 00655: MOV_11
    "10000011",
    "00001000",  -- 00657: INC_2
    "10000110",  -- 00658: MOV_11
    "11110000",
    "00001000",  -- 00660: INC_2
    "11100110",  -- 00661: MOV_3
    "00010010",  -- 00662: LCALL
    "00000011",
    "01000011",
    "10101100",  -- 00665: MOV_6
    "10000010",
    "10101101",  -- 00667: MOV_6
    "10000011",
    "10101110",  -- 00669: MOV_6
    "11110000",
    "11111111",  -- 00671: MOV_5
    "11100101",  -- 00672: MOV_2
    "10000001",
    "00100100",  -- 00674: ADD_4
    "11111100",
    "11110101",  -- 00676: MOV_8
    "10000001",
    "11100101",  -- 00678: MOV_2
    "00001000",
    "00100100",  -- 00680: ADD_4
    "00001001",
    "11111000",  -- 00682: MOV_5
    "11100110",  -- 00683: MOV_3
    "00110000",  -- 00684: JNB
    "11100000",
    "00101011",
    "11000000",  -- 00687: PUSH
    "00000100",
    "11000000",  -- 00689: PUSH
    "00000101",
    "11000000",  -- 00691: PUSH
    "00000110",
    "11000000",  -- 00693: PUSH
    "00000111",
    "10010000",  -- 00695: MOV_18
    "00000100",
    "11110011",
    "01110101",  -- 00698: MOV_12
    "11110000",
    "00110101",
    "01110100",  -- 00701: MOV_4
    "00111111",
    "00010010",  -- 00703: LCALL
    "00000110",
    "10100011",
    "10101100",  -- 00706: MOV_6
    "10000010",
    "10101101",  -- 00708: MOV_6
    "10000011",
    "10101110",  -- 00710: MOV_6
    "11110000",
    "11111111",  -- 00712: MOV_5
    "11100101",  -- 00713: MOV_2
    "10000001",
    "00100100",  -- 00715: ADD_4
    "11111100",
    "11110101",  -- 00717: MOV_8
    "10000001",
    "11100101",  -- 00719: MOV_2
    "00001000",
    "00100100",  -- 00721: ADD_4
    "00001001",
    "11111000",  -- 00723: MOV_5
    "00000110",  -- 00724: INC_4
    "10110110",  -- 00725: CJNE_4
    "00000000",
    "00000010",
    "00001000",  -- 00728: INC_2
    "00000110",  -- 00729: INC_4
    "01110101",  -- 00730: MOV_12
    "00001011",
    "00000010",
    "01110101",  -- 00733: MOV_12
    "00001100",
    "00000000",
    "11100101",  -- 00736: MOV_2
    "00001000",
    "00100100",  -- 00738: ADD_4
    "00001001",
    "11111000",  -- 00740: MOV_5
    "10000110",  -- 00741: MOV_11
    "10000010",
    "00001000",  -- 00743: INC_2
    "10000110",  -- 00744: MOV_11
    "10000011",
    "11000000",  -- 00746: PUSH
    "00000111",
    "11000000",  -- 00748: PUSH
    "00000110",
    "11000000",  -- 00750: PUSH
    "00000101",
    "11000000",  -- 00752: PUSH
    "00000100",
    "00010010",  -- 00754: LCALL
    "00000110",
    "01101011",
    "10000101",  -- 00757: MOV_10
    "10000010",
    "00001011",
    "10000101",  -- 00760: MOV_10
    "10000011",
    "00001100",
    "11010000",  -- 00763: POP
    "00000100",
    "11010000",  -- 00765: POP
    "00000101",
    "11010000",  -- 00767: POP
    "00000110",
    "11010000",  -- 00769: POP
    "00000111",
    "10001100",  -- 00771: MOV_9
    "10000010",
    "10001101",  -- 00773: MOV_9
    "10000011",
    "10001110",  -- 00775: MOV_9
    "11110000",
    "11101111",  -- 00777: MOV_1
    "00010010",  -- 00778: LCALL
    "00000011",
    "11000101",
    "10000101",  -- 00781: MOV_10
    "00001000",
    "10000001",
    "11010000",  -- 00784: POP
    "00001000",
    "00100010",  -- 00786: RET
    "11111111",  -- 00787: MOV_5
    "10101000",  -- 00788: MOV_6
    "10000001",
    "00011000",  -- 00790: DEC_2
    "00011000",  -- 00791: DEC_2
    "00010010",  -- 00792: LCALL
    "00000100",
    "01110111",
    "11010010",  -- 00795: SETB_2
    "11010001",
    "00110011",  -- 00797: RLC
    "11100110",  -- 00798: MOV_3
    "01000000",  -- 00799: JC
    "00000111",
    "00110000",  -- 00801: JNB
    "11100111",
    "00001011",
    "01110101",  -- 00804: MOV_12
    "10000010",
    "00000000",
    "00100010",  -- 00807: RET
    "00100000",  -- 00808: JB
    "11100111",
    "00000110",
    "01110101",  -- 00811: MOV_12
    "10000010",
    "00000001",
    "00100010",  -- 00814: RET
    "11000010",  -- 00815: CLR_3
    "11010001",
    "00010010",  -- 00817: LCALL
    "00000100",
    "01011001",
    "11101001",  -- 00820: MOV_1
    "01110000",  -- 00821: JNZ
    "00000011",
    "11110101",  -- 00823: MOV_8
    "10000010",
    "00100010",  -- 00825: RET
    "00100000",  -- 00826: JB
    "11010001",
    "00000001",
    "10110011",  -- 00829: CPL_2
    "11100100",  -- 00830: CLR_1
    "00110011",  -- 00831: RLC
    "11110101",  -- 00832: MOV_8
    "10000010",
    "00100010",  -- 00834: RET
    "00010010",  -- 00835: LCALL
    "00000111",
    "01000110",
    "01111001",  -- 00838: MOV_7
    "00000000",
    "11100101",  -- 00840: MOV_2
    "10000011",
    "10110101",  -- 00842: CJNE_1
    "10000010",
    "00000010",
    "10000000",  -- 00845: SJMP
    "00001101",
    "01010000",  -- 00847: JNC
    "00000011",
    "00010010",  -- 00849: LCALL
    "00000101",
    "10000110",
    "11100101",  -- 00852: MOV_2
    "10000011",
    "11000011",  -- 00854: CLR_2
    "10010101",  -- 00855: SUBB_2
    "10000010",
    "00010010",  -- 00857: LCALL
    "00000111",
    "01110100",
    "11100101",  -- 00860: MOV_2
    "11010000",
    "11000100",  -- 00862: SWAP
    "01100101",  -- 00863: XRL_2
    "11010000",
    "00100000",  -- 00865: JB
    "11100001",
    "00010111",
    "11101010",  -- 00868: MOV_1
    "00101101",  -- 00869: ADD_1
    "11111010",  -- 00870: MOV_5
    "11101011",  -- 00871: MOV_1
    "00111110",  -- 00872: ADDC_1
    "11111011",  -- 00873: MOV_5
    "11101100",  -- 00874: MOV_1
    "00111111",  -- 00875: ADDC_1
    "11111100",  -- 00876: MOV_5
    "01010000",  -- 00877: JNC
    "00001001",
    "01110100",  -- 00879: MOV_4
    "00000001",
    "00010010",  -- 00881: LCALL
    "00000111",
    "01110100",
    "11101100",  -- 00884: MOV_1
    "01000100",  -- 00885: ORL_4
    "10000000",
    "11111100",  -- 00887: MOV_5
    "00000010",  -- 00888: LJMP
    "00000101",
    "00110111",
    "11000011",  -- 00891: CLR_2
    "11101010",  -- 00892: MOV_1
    "10011101",  -- 00893: SUBB_1
    "11111010",  -- 00894: MOV_5
    "11101011",  -- 00895: MOV_1
    "10011110",  -- 00896: SUBB_1
    "11111011",  -- 00897: MOV_5
    "11101100",  -- 00898: MOV_1
    "10011111",  -- 00899: SUBB_1
    "11111100",  -- 00900: MOV_5
    "01010000",  -- 00901: JNC
    "00001111",
    "11000011",  -- 00903: CLR_2
    "11100100",  -- 00904: CLR_1
    "10011001",  -- 00905: SUBB_1
    "11111001",  -- 00906: MOV_5
    "11100100",  -- 00907: CLR_1
    "10011010",  -- 00908: SUBB_1
    "11111010",  -- 00909: MOV_5
    "11100100",  -- 00910: CLR_1
    "10011011",  -- 00911: SUBB_1
    "11111011",  -- 00912: MOV_5
    "11100100",  -- 00913: CLR_1
    "10011100",  -- 00914: SUBB_1
    "11111100",  -- 00915: MOV_5
    "10110010",  -- 00916: CPL_3
    "11010001",
    "00010010",  -- 00918: LCALL
    "00000111",
    "10110111",
    "00000010",  -- 00921: LJMP
    "00000101",
    "00110111",
    "01111010",  -- 00924: MOV_7
    "00010000",
    "11100100",  -- 00926: CLR_1
    "11111011",  -- 00927: MOV_5
    "11111100",  -- 00928: MOV_5
    "11100101",  -- 00929: MOV_2
    "10000010",
    "00100101",  -- 00931: ADD_2
    "11100000",
    "11110101",  -- 00933: MOV_8
    "10000010",
    "11100101",  -- 00935: MOV_2
    "10000011",
    "00110011",  -- 00937: RLC
    "11110101",  -- 00938: MOV_8
    "10000011",
    "11101011",  -- 00940: MOV_1
    "00110011",  -- 00941: RLC
    "11111011",  -- 00942: MOV_5
    "11101100",  -- 00943: MOV_1
    "00110011",  -- 00944: RLC
    "11111100",  -- 00945: MOV_5
    "11101011",  -- 00946: MOV_1
    "10010101",  -- 00947: SUBB_2
    "00001011",
    "11110101",  -- 00949: MOV_8
    "11110000",
    "11101100",  -- 00951: MOV_1
    "10010101",  -- 00952: SUBB_2
    "00001100",
    "01000000",  -- 00954: JC
    "00000110",
    "11111100",  -- 00956: MOV_5
    "10101011",  -- 00957: MOV_6
    "11110000",
    "01000011",  -- 00959: ORL_6
    "10000010",
    "00000001",
    "11011010",  -- 00962: DJNZ_1
    "11011101",
    "00100010",  -- 00964: RET
    "10101100",  -- 00965: MOV_6
    "10000010",
    "10101101",  -- 00967: MOV_6
    "10000011",
    "10101110",  -- 00969: MOV_6
    "11110000",
    "11111111",  -- 00971: MOV_5
    "10001100",  -- 00972: MOV_9
    "00001101",
    "10001101",  -- 00974: MOV_9
    "00001110",
    "10001110",  -- 00976: MOV_9
    "00001111",
    "10001111",  -- 00978: MOV_9
    "00010000",
    "10101100",  -- 00980: MOV_6
    "00001101",
    "10101101",  -- 00982: MOV_6
    "00001110",
    "10101110",  -- 00984: MOV_6
    "00001111",
    "10101111",  -- 00986: MOV_6
    "00010000",
    "10001110",  -- 00988: MOV_9
    "00000100",
    "11101111",  -- 00990: MOV_1
    "10100010",  -- 00991: MOV_16
    "11100111",
    "11001100",  -- 00993: XCH_1
    "00110011",  -- 00994: RLC
    "11001100",  -- 00995: XCH_1
    "00110011",  -- 00996: RLC
    "11001100",  -- 00997: XCH_1
    "01010100",  -- 00998: ANL_4
    "00000001",
    "00110000",  -- 01000: JNB
    "11100000",
    "00000010",
    "01000100",  -- 01003: ORL_4
    "11111110",
    "00110011",  -- 01005: RLC
    "10010101",  -- 01006: SUBB_2
    "11100000",
    "10001100",  -- 01008: MOV_9
    "00010001",
    "01110101",  -- 01010: MOV_12
    "00010010",
    "00000000",
    "01110101",  -- 01013: MOV_12
    "00010011",
    "00000000",
    "01110101",  -- 01016: MOV_12
    "00010100",
    "00000000",
    "10101010",  -- 01019: MOV_6
    "00001011",
    "11100101",  -- 01021: MOV_2
    "00001100",
    "11111011",  -- 01023: MOV_5
    "00110011",  -- 01024: RLC
    "10010101",  -- 01025: SUBB_2
    "11100000",
    "11111110",  -- 01027: MOV_5
    "11111111",  -- 01028: MOV_5
    "11101010",  -- 01029: MOV_1
    "00100101",  -- 01030: ADD_2
    "00010001",
    "11111010",  -- 01032: MOV_5
    "11101011",  -- 01033: MOV_1
    "00110101",  -- 01034: ADDC_2
    "00010010",
    "11101110",  -- 01036: MOV_1
    "00110101",  -- 01037: ADDC_2
    "00010011",
    "11101111",  -- 01039: MOV_1
    "00110101",  -- 01040: ADDC_2
    "00010100",
    "01111011",  -- 01042: MOV_7
    "00000000",
    "10001010",  -- 01044: MOV_9
    "00010011",
    "11101011",  -- 01046: MOV_1
    "01010100",  -- 01047: ANL_4
    "00000001",
    "10100010",  -- 01049: MOV_16
    "11100000",
    "11000101",  -- 01051: XCH_2
    "00010011",
    "00010011",  -- 01053: RRC
    "11000101",  -- 01054: XCH_2
    "00010011",
    "00010011",  -- 01056: RRC
    "11000101",  -- 01057: XCH_2
    "00010011",
    "11110101",  -- 01059: MOV_8
    "00010100",
    "01110101",  -- 01061: MOV_12
    "00010001",
    "00000000",
    "01110101",  -- 01064: MOV_12
    "00010010",
    "00000000",
    "10101100",  -- 01067: MOV_6
    "00001101",
    "10101101",  -- 01069: MOV_6
    "00001110",
    "10101110",  -- 01071: MOV_6
    "00001111",
    "10101111",  -- 01073: MOV_6
    "00010000",
    "01010011",  -- 01075: ANL_6
    "00000110",
    "01111111",
    "01010011",  -- 01078: ANL_6
    "00000111",
    "10000000",
    "11100101",  -- 01081: MOV_2
    "00010011",
    "01000010",  -- 01083: ORL_5
    "00000110",
    "11100101",  -- 01085: MOV_2
    "00010100",
    "01000010",  -- 01087: ORL_5
    "00000111",
    "10001100",  -- 01089: MOV_9
    "00001101",
    "10001101",  -- 01091: MOV_9
    "00001110",
    "10001110",  -- 01093: MOV_9
    "00001111",
    "10001111",  -- 01095: MOV_9
    "00010000",
    "10101100",  -- 01097: MOV_6
    "00001101",
    "10101101",  -- 01099: MOV_6
    "00001110",
    "10101110",  -- 01101: MOV_6
    "00001111",
    "10101111",  -- 01103: MOV_6
    "00010000",
    "10001100",  -- 01105: MOV_9
    "10000010",
    "10001101",  -- 01107: MOV_9
    "10000011",
    "10001110",  -- 01109: MOV_9
    "11110000",
    "11101111",  -- 01111: MOV_1
    "00100010",  -- 01112: RET
    "01111001",  -- 01113: MOV_7
    "00000001",
    "10101010",  -- 01115: MOV_6
    "10000010",
    "11100110",  -- 01117: MOV_3
    "10001111",  -- 01118: MOV_9
    "10000010",
    "10110101",  -- 01120: CJNE_1
    "10000010",
    "00010011",
    "00011000",  -- 01123: DEC_2
    "11100110",  -- 01124: MOV_3
    "10110101",  -- 01125: CJNE_1
    "11110000",
    "00001110",
    "00011000",  -- 01128: DEC_2
    "11100110",  -- 01129: MOV_3
    "10110101",  -- 01130: CJNE_1
    "10000011",
    "00001001",
    "00011000",  -- 01133: DEC_2
    "11100110",  -- 01134: MOV_3
    "10001010",  -- 01135: MOV_9
    "10000010",
    "10110101",  -- 01137: CJNE_1
    "10000010",
    "00000010",
    "01111001",  -- 01140: MOV_7
    "00000000",
    "00100010",  -- 01142: RET
    "10110100",  -- 01143: CJNE_2
    "10000000",
    "00001111",
    "11100101",  -- 01146: MOV_2
    "11110000",
    "01110000",  -- 01148: JNZ
    "00001010",
    "11100101",  -- 01150: MOV_2
    "10000011",
    "01110000",  -- 01152: JNZ
    "00000110",
    "11100101",  -- 01154: MOV_2
    "10000010",
    "01110000",  -- 01156: JNZ
    "00000010",
    "01111111",  -- 01158: MOV_7
    "00000000",
    "11101111",  -- 01160: MOV_1
    "10110110",  -- 01161: CJNE_4
    "10000000",
    "00010101",
    "00011000",  -- 01164: DEC_2
    "10110110",  -- 01165: CJNE_4
    "00000000",
    "00010000",
    "00011000",  -- 01168: DEC_2
    "10110110",  -- 01169: CJNE_4
    "00000000",
    "00001011",
    "00011000",  -- 01172: DEC_2
    "10110110",  -- 01173: CJNE_4
    "00000000",
    "00000110",
    "00001000",  -- 01176: INC_2
    "00001000",  -- 01177: INC_2
    "00001000",  -- 01178: INC_2
    "01110110",  -- 01179: MOV_15
    "00000000",
    "00100010",  -- 01181: RET
    "00001000",  -- 01182: INC_2
    "00001000",  -- 01183: INC_2
    "00001000",  -- 01184: INC_2
    "00100010",  -- 01185: RET
    "10101100",  -- 01186: MOV_6
    "10000010",
    "10101101",  -- 01188: MOV_6
    "10000011",
    "10101110",  -- 01190: MOV_6
    "11110000",
    "11111111",  -- 01192: MOV_5
    "10001100",  -- 01193: MOV_9
    "00001110",
    "10001101",  -- 01195: MOV_9
    "00001111",
    "10001110",  -- 01197: MOV_9
    "00010000",
    "10001111",  -- 01199: MOV_9
    "00010001",
    "10101100",  -- 01201: MOV_6
    "00001110",
    "10101101",  -- 01203: MOV_6
    "00001111",
    "10101110",  -- 01205: MOV_6
    "00010000",
    "10101111",  -- 01207: MOV_6
    "00010001",
    "10001110",  -- 01209: MOV_9
    "00000100",
    "11101111",  -- 01211: MOV_1
    "10100010",  -- 01212: MOV_16
    "11100111",
    "11001100",  -- 01214: XCH_1
    "00110011",  -- 01215: RLC
    "11001100",  -- 01216: XCH_1
    "00110011",  -- 01217: RLC
    "11001100",  -- 01218: XCH_1
    "01010100",  -- 01219: ANL_4
    "00000001",
    "00110000",  -- 01221: JNB
    "11100000",
    "00000010",
    "01000100",  -- 01224: ORL_4
    "11111110",
    "00110011",  -- 01226: RLC
    "10010101",  -- 01227: SUBB_2
    "11100000",
    "11100100",  -- 01229: CLR_1
    "11111101",  -- 01230: MOV_5
    "11111110",  -- 01231: MOV_5
    "11111111",  -- 01232: MOV_5
    "11101100",  -- 01233: MOV_1
    "00100100",  -- 01234: ADD_4
    "10000010",
    "11110101",  -- 01236: MOV_8
    "00010010",
    "11101101",  -- 01238: MOV_1
    "00110100",  -- 01239: ADDC_4
    "11111111",
    "11110101",  -- 01241: MOV_8
    "00010011",
    "11101110",  -- 01243: MOV_1
    "00110100",  -- 01244: ADDC_4
    "11111111",
    "11110101",  -- 01246: MOV_8
    "00010100",
    "11101111",  -- 01248: MOV_1
    "00110100",  -- 01249: ADDC_4
    "11111111",
    "11110101",  -- 01251: MOV_8
    "00010101",
    "10101010",  -- 01253: MOV_6
    "00001011",
    "10101011",  -- 01255: MOV_6
    "00001100",
    "10101111",  -- 01257: MOV_6
    "00001101",
    "10101100",  -- 01259: MOV_6
    "00010010",
    "10101101",  -- 01261: MOV_6
    "00010011",
    "10001010",  -- 01263: MOV_9
    "10000010",
    "10001011",  -- 01265: MOV_9
    "10000011",
    "10001111",  -- 01267: MOV_9
    "11110000",
    "11101100",  -- 01269: MOV_1
    "00010010",  -- 01270: LCALL
    "00001000",
    "00100010",
    "10100011",  -- 01273: INC_5
    "11101101",  -- 01274: MOV_1
    "00010010",  -- 01275: LCALL
    "00001000",
    "00100010",
    "10101100",  -- 01278: MOV_6
    "00001110",
    "10101101",  -- 01280: MOV_6
    "00001111",
    "10101110",  -- 01282: MOV_6
    "00010000",
    "10101111",  -- 01284: MOV_6
    "00010001",
    "01010011",  -- 01286: ANL_6
    "00000110",
    "01111111",
    "01010011",  -- 01289: ANL_6
    "00000111",
    "10000000",
    "10001100",  -- 01292: MOV_9
    "00001110",
    "10001101",  -- 01294: MOV_9
    "00001111",
    "10001110",  -- 01296: MOV_9
    "00010000",
    "10001111",  -- 01298: MOV_9
    "00010001",
    "10101100",  -- 01300: MOV_6
    "00001110",
    "10101101",  -- 01302: MOV_6
    "00001111",
    "10101110",  -- 01304: MOV_6
    "00010000",
    "10101111",  -- 01306: MOV_6
    "00010001",
    "01000011",  -- 01308: ORL_6
    "00000111",
    "00111111",
    "10001100",  -- 01311: MOV_9
    "00001110",
    "10001101",  -- 01313: MOV_9
    "00001111",
    "10001110",  -- 01315: MOV_9
    "00010000",
    "10001111",  -- 01317: MOV_9
    "00010001",
    "10101100",  -- 01319: MOV_6
    "00001110",
    "10101101",  -- 01321: MOV_6
    "00001111",
    "10101110",  -- 01323: MOV_6
    "00010000",
    "10101111",  -- 01325: MOV_6
    "00010001",
    "10001100",  -- 01327: MOV_9
    "10000010",
    "10001101",  -- 01329: MOV_9
    "10000011",
    "10001110",  -- 01331: MOV_9
    "11110000",
    "11101111",  -- 01333: MOV_1
    "00100010",  -- 01334: RET
    "10111001",  -- 01335: CJNE_3
    "10000000",
    "00000011",
    "11101010",  -- 01338: MOV_1
    "00010011",  -- 01339: RRC
    "10110011",  -- 01340: CPL_2
    "01000000",  -- 01341: JC
    "00010000",
    "11101010",  -- 01343: MOV_1
    "00100100",  -- 01344: ADD_4
    "00000001",
    "11111010",  -- 01346: MOV_5
    "11100100",  -- 01347: CLR_1
    "00111011",  -- 01348: ADDC_1
    "11111011",  -- 01349: MOV_5
    "11100100",  -- 01350: CLR_1
    "00111100",  -- 01351: ADDC_1
    "11111100",  -- 01352: MOV_5
    "01010000",  -- 01353: JNC
    "00000100",
    "01111100",  -- 01355: MOV_7
    "10000000",
    "00000101",  -- 01357: INC_3
    "10000010",
    "10111100",  -- 01359: CJNE_3
    "00000000",
    "00001110",
    "10111011",  -- 01362: CJNE_3
    "00000000",
    "00001011",
    "10111010",  -- 01365: CJNE_3
    "00000000",
    "00001000",
    "11100100",  -- 01368: CLR_1
    "11110101",  -- 01369: MOV_8
    "11110000",
    "11110101",  -- 01371: MOV_8
    "10000011",
    "11110101",  -- 01373: MOV_8
    "10000010",
    "00100010",  -- 01375: RET
    "10100010",  -- 01376: MOV_16
    "11010001",
    "11100101",  -- 01378: MOV_2
    "10000010",
    "00010011",  -- 01380: RRC
    "10001100",  -- 01381: MOV_9
    "11110000",
    "10010010",  -- 01383: MOV_17
    "11110111",
    "10001011",  -- 01385: MOV_9
    "10000011",
    "10001010",  -- 01387: MOV_9
    "10000010",
    "00100010",  -- 01389: RET
    "11100100",  -- 01390: CLR_1
    "11110101",  -- 01391: MOV_8
    "10000011",
    "11110101",  -- 01393: MOV_8
    "10000010",
    "01110101",  -- 01395: MOV_12
    "11110000",
    "10000000",
    "11110100",  -- 01398: CPL_1
    "10100010",  -- 01399: MOV_16
    "11010001",
    "00010011",  -- 01401: RRC
    "00100010",  -- 01402: RET
    "11100100",  -- 01403: CLR_1
    "11110101",  -- 01404: MOV_8
    "10000011",
    "11110101",  -- 01406: MOV_8
    "10000010",
    "01110101",  -- 01408: MOV_12
    "11110000",
    "11000000",
    "01110100",  -- 01411: MOV_4
    "01111111",
    "00100010",  -- 01413: RET
    "11100101",  -- 01414: MOV_2
    "10000010",
    "11000101",  -- 01416: XCH_2
    "10000011",
    "11110101",  -- 01418: MOV_8
    "10000010",
    "10100010",  -- 01420: MOV_16
    "11010001",
    "00110011",  -- 01422: RLC
    "10100010",  -- 01423: MOV_16
    "11010101",
    "10010010",  -- 01425: MOV_17
    "11010001",
    "00010011",  -- 01427: RRC
    "10010010",  -- 01428: MOV_17
    "11010101",
    "11101100",  -- 01430: MOV_1
    "11001111",  -- 01431: XCH_1
    "11111100",  -- 01432: MOV_5
    "11101011",  -- 01433: MOV_1
    "11001110",  -- 01434: XCH_1
    "11111011",  -- 01435: MOV_5
    "11101010",  -- 01436: MOV_1
    "11001101",  -- 01437: XCH_1
    "11111010",  -- 01438: MOV_5
    "00100010",  -- 01439: RET
    "00010010",  -- 01440: LCALL
    "00000111",
    "01000110",
    "00110000",  -- 01443: JNB
    "11010101",
    "00000010",
    "10110010",  -- 01446: CPL_3
    "11010001",
    "10111111",  -- 01448: CJNE_3
    "00000000",
    "00001001",
    "10111100",  -- 01451: CJNE_3
    "00000000",
    "00000011",
    "00000010",  -- 01454: LJMP
    "00000101",
    "01111011",
    "00000010",  -- 01457: LJMP
    "00000101",
    "01101110",
    "10111100",  -- 01460: CJNE_3
    "00000000",
    "00000011",
    "00000010",  -- 01463: LJMP
    "00000101",
    "01011000",
    "11100101",  -- 01466: MOV_2
    "10000011",
    "10110100",  -- 01468: CJNE_2
    "11111111",
    "00001011",
    "11100101",  -- 01471: MOV_2
    "10000010",
    "10110100",  -- 01473: CJNE_2
    "11111111",
    "00000011",
    "00000010",  -- 01476: LJMP
    "00000101",
    "01111011",
    "00000010",  -- 01479: LJMP
    "00000101",
    "01011000",
    "11100101",  -- 01482: MOV_2
    "10000010",
    "10110100",  -- 01484: CJNE_2
    "11111111",
    "00000011",
    "00000010",  -- 01487: LJMP
    "00000101",
    "01101110",
    "11000011",  -- 01490: CLR_2
    "10010101",  -- 01491: SUBB_2
    "10000011",
    "01010000",  -- 01493: JNC
    "00000111",
    "00100100",  -- 01495: ADD_4
    "01111111",
    "01000000",  -- 01497: JC
    "00001011",
    "00000010",  -- 01499: LJMP
    "00000101",
    "01011000",
    "00100100",  -- 01502: ADD_4
    "10000000",
    "00010100",  -- 01504: DEC_1
    "01010000",  -- 01505: JNC
    "00000011",
    "00000010",  -- 01507: LJMP
    "00000101",
    "01101110",
    "11110101",  -- 01510: MOV_8
    "10000010",
    "11000011",  -- 01512: CLR_2
    "11101101",  -- 01513: MOV_1
    "10011010",  -- 01514: SUBB_1
    "11101110",  -- 01515: MOV_1
    "10011011",  -- 01516: SUBB_1
    "11101111",  -- 01517: MOV_1
    "10011100",  -- 01518: SUBB_1
    "01000000",  -- 01519: JC
    "00010001",
    "00010101",  -- 01521: DEC_3
    "10000010",
    "11000011",  -- 01523: CLR_2
    "11101010",  -- 01524: MOV_1
    "00110011",  -- 01525: RLC
    "11111001",  -- 01526: MOV_5
    "11101011",  -- 01527: MOV_1
    "00110011",  -- 01528: RLC
    "11111010",  -- 01529: MOV_5
    "11101100",  -- 01530: MOV_1
    "00110011",  -- 01531: RLC
    "11111011",  -- 01532: MOV_5
    "11100100",  -- 01533: CLR_1
    "00110011",  -- 01534: RLC
    "11111100",  -- 01535: MOV_5
    "10000000",  -- 01536: SJMP
    "00000101",
    "11100100",  -- 01538: CLR_1
    "11001100",  -- 01539: XCH_1
    "11001011",  -- 01540: XCH_1
    "11001010",  -- 01541: XCH_1
    "11111001",  -- 01542: MOV_5
    "11000000",  -- 01543: PUSH
    "10000010",
    "01110101",  -- 01545: MOV_12
    "11110000",
    "00011001",
    "11000011",  -- 01548: CLR_2
    "11101001",  -- 01549: MOV_1
    "10011101",  -- 01550: SUBB_1
    "11101010",  -- 01551: MOV_1
    "10011110",  -- 01552: SUBB_1
    "11101011",  -- 01553: MOV_1
    "10011111",  -- 01554: SUBB_1
    "11101100",  -- 01555: MOV_1
    "10010100",  -- 01556: SUBB_4
    "00000000",
    "11010101",  -- 01558: DJNZ_2
    "11110000",
    "00000010",
    "10000000",  -- 01561: SJMP
    "00101101",
    "01000000",  -- 01563: JC
    "00001110",
    "11101001",  -- 01565: MOV_1
    "10011101",  -- 01566: SUBB_1
    "11111001",  -- 01567: MOV_5
    "11101010",  -- 01568: MOV_1
    "10011110",  -- 01569: SUBB_1
    "11111010",  -- 01570: MOV_5
    "11101011",  -- 01571: MOV_1
    "10011111",  -- 01572: SUBB_1
    "11111011",  -- 01573: MOV_5
    "11101100",  -- 01574: MOV_1
    "10010100",  -- 01575: SUBB_4
    "00000000",
    "11111100",  -- 01577: MOV_5
    "11000011",  -- 01578: CLR_2
    "10110011",  -- 01579: CPL_2
    "11101000",  -- 01580: MOV_1
    "00110011",  -- 01581: RLC
    "11111000",  -- 01582: MOV_5
    "11100101",  -- 01583: MOV_2
    "10000010",
    "00110011",  -- 01585: RLC
    "11110101",  -- 01586: MOV_8
    "10000010",
    "11100101",  -- 01588: MOV_2
    "10000011",
    "00110011",  -- 01590: RLC
    "11110101",  -- 01591: MOV_8
    "10000011",
    "11000011",  -- 01593: CLR_2
    "11101001",  -- 01594: MOV_1
    "00110011",  -- 01595: RLC
    "11111001",  -- 01596: MOV_5
    "11101010",  -- 01597: MOV_1
    "00110011",  -- 01598: RLC
    "11111010",  -- 01599: MOV_5
    "11101011",  -- 01600: MOV_1
    "00110011",  -- 01601: RLC
    "11111011",  -- 01602: MOV_5
    "11101100",  -- 01603: MOV_1
    "00110011",  -- 01604: RLC
    "11111100",  -- 01605: MOV_5
    "10000000",  -- 01606: SJMP
    "11000100",
    "10110011",  -- 01608: CPL_2
    "11100100",  -- 01609: CLR_1
    "11111001",  -- 01610: MOV_5
    "00111000",  -- 01611: ADDC_1
    "11111010",  -- 01612: MOV_5
    "11100100",  -- 01613: CLR_1
    "00110101",  -- 01614: ADDC_2
    "10000010",
    "11111011",  -- 01616: MOV_5
    "11100100",  -- 01617: CLR_1
    "00110101",  -- 01618: ADDC_2
    "10000011",
    "11111100",  -- 01620: MOV_5
    "11010000",  -- 01621: POP
    "10000010",
    "01010000",  -- 01623: JNC
    "00000100",
    "00000101",  -- 01625: INC_3
    "10000010",
    "01111100",  -- 01627: MOV_7
    "10000000",
    "00010010",  -- 01629: LCALL
    "00000111",
    "10110111",
    "00000010",  -- 01632: LJMP
    "00000101",
    "01001111",
    "01111111",  -- 01635: MOV_7
    "10000110",
    "00010010",  -- 01637: LCALL
    "00000111",
    "11111101",
    "11110101",  -- 01640: MOV_8
    "10000010",
    "00100010",  -- 01642: RET
    "11000010",  -- 01643: CLR_3
    "11010101",
    "11100101",  -- 01645: MOV_2
    "10000011",
    "00110000",  -- 01647: JNB
    "11100111",
    "00001101",
    "11010010",  -- 01650: SETB_2
    "11010101",
    "11100100",  -- 01652: CLR_1
    "11000011",  -- 01653: CLR_2
    "10010101",  -- 01654: SUBB_2
    "10000010",
    "11110101",  -- 01656: MOV_8
    "10000010",
    "11100100",  -- 01658: CLR_1
    "10010101",  -- 01659: SUBB_2
    "10000011",
    "11110101",  -- 01661: MOV_8
    "10000011",
    "11100101",  -- 01663: MOV_2
    "00001100",
    "00110000",  -- 01665: JNB
    "11100111",
    "00001101",
    "10110010",  -- 01668: CPL_3
    "11010101",
    "11100100",  -- 01670: CLR_1
    "11000011",  -- 01671: CLR_2
    "10010101",  -- 01672: SUBB_2
    "00001011",
    "11110101",  -- 01674: MOV_8
    "00001011",
    "11100100",  -- 01676: CLR_1
    "10010101",  -- 01677: SUBB_2
    "00001100",
    "11110101",  -- 01679: MOV_8
    "00001100",
    "00010010",  -- 01681: LCALL
    "00000011",
    "10011100",
    "00110000",  -- 01684: JNB
    "11010101",
    "00001011",
    "11100100",  -- 01687: CLR_1
    "11000011",  -- 01688: CLR_2
    "10010101",  -- 01689: SUBB_2
    "10000010",
    "11110101",  -- 01691: MOV_8
    "10000010",
    "11100100",  -- 01693: CLR_1
    "10010101",  -- 01694: SUBB_2
    "10000011",
    "11110101",  -- 01696: MOV_8
    "10000011",
    "00100010",  -- 01698: RET
    "00010010",  -- 01699: LCALL
    "00000111",
    "01000110",
    "10111100",  -- 01702: CJNE_3
    "00000000",
    "00000011",
    "00000010",  -- 01705: LJMP
    "00000101",
    "01011000",
    "11101111",  -- 01708: MOV_1
    "01100000",  -- 01709: JZ
    "11111010",
    "00110000",  -- 01711: JNB
    "11010101",
    "00000010",
    "10110010",  -- 01714: CPL_3
    "11010001",
    "11100101",  -- 01716: MOV_2
    "10000011",
    "10110100",  -- 01718: CJNE_2
    "11111111",
    "00000011",
    "00000010",  -- 01721: LJMP
    "00000101",
    "01101110",
    "11100101",  -- 01724: MOV_2
    "10000010",
    "10110100",  -- 01726: CJNE_2
    "11111111",
    "00000011",
    "00000010",  -- 01729: LJMP
    "00000101",
    "01101110",
    "00100101",  -- 01732: ADD_2
    "10000011",
    "01000000",  -- 01734: JC
    "00000111",
    "00100100",  -- 01736: ADD_4
    "10000010",
    "01000000",  -- 01738: JC
    "00001011",
    "00000010",  -- 01740: LJMP
    "00000101",
    "01011000",
    "00100100",  -- 01743: ADD_4
    "10000011",
    "00010100",  -- 01745: DEC_1
    "01010000",  -- 01746: JNC
    "00000011",
    "00000010",  -- 01748: LJMP
    "00000101",
    "01101110",
    "11110101",  -- 01751: MOV_8
    "10000010",
    "11101010",  -- 01753: MOV_1
    "10001101",  -- 01754: MOV_9
    "11110000",
    "10100100",  -- 01756: MUL
    "10101000",  -- 01757: MOV_6
    "11110000",
    "11101010",  -- 01759: MOV_1
    "10001110",  -- 01760: MOV_9
    "11110000",
    "10100100",  -- 01762: MUL
    "00101000",  -- 01763: ADD_1
    "11111000",  -- 01764: MOV_5
    "11100100",  -- 01765: CLR_1
    "00110101",  -- 01766: ADDC_2
    "11110000",
    "11111001",  -- 01768: MOV_5
    "11101011",  -- 01769: MOV_1
    "10001101",  -- 01770: MOV_9
    "11110000",
    "10100100",  -- 01772: MUL
    "00101000",  -- 01773: ADD_1
    "11101001",  -- 01774: MOV_1
    "00110101",  -- 01775: ADDC_2
    "11110000",
    "11111001",  -- 01777: MOV_5
    "11100100",  -- 01778: CLR_1
    "00110011",  -- 01779: RLC
    "11001010",  -- 01780: XCH_1
    "10001111",  -- 01781: MOV_9
    "11110000",
    "10100100",  -- 01783: MUL
    "00101001",  -- 01784: ADD_1
    "11111001",  -- 01785: MOV_5
    "11101010",  -- 01786: MOV_1
    "00110101",  -- 01787: ADDC_2
    "11110000",
    "11111010",  -- 01789: MOV_5
    "11101011",  -- 01790: MOV_1
    "11111000",  -- 01791: MOV_5
    "10001110",  -- 01792: MOV_9
    "11110000",
    "10100100",  -- 01794: MUL
    "00101001",  -- 01795: ADD_1
    "11111001",  -- 01796: MOV_5
    "11101010",  -- 01797: MOV_1
    "00110101",  -- 01798: ADDC_2
    "11110000",
    "11111010",  -- 01800: MOV_5
    "11100100",  -- 01801: CLR_1
    "00110011",  -- 01802: RLC
    "11111011",  -- 01803: MOV_5
    "11101100",  -- 01804: MOV_1
    "10001101",  -- 01805: MOV_9
    "11110000",
    "10100100",  -- 01807: MUL
    "00101001",  -- 01808: ADD_1
    "11111001",  -- 01809: MOV_5
    "11101010",  -- 01810: MOV_1
    "00110101",  -- 01811: ADDC_2
    "11110000",
    "11111010",  -- 01813: MOV_5
    "11100100",  -- 01814: CLR_1
    "00111011",  -- 01815: ADDC_1
    "11111011",  -- 01816: MOV_5
    "11101000",  -- 01817: MOV_1
    "10001111",  -- 01818: MOV_9
    "11110000",
    "10100100",  -- 01820: MUL
    "00101010",  -- 01821: ADD_1
    "11111010",  -- 01822: MOV_5
    "11101011",  -- 01823: MOV_1
    "00110101",  -- 01824: ADDC_2
    "11110000",
    "11111011",  -- 01826: MOV_5
    "11100100",  -- 01827: CLR_1
    "00110011",  -- 01828: RLC
    "11001100",  -- 01829: XCH_1
    "11111101",  -- 01830: MOV_5
    "10001110",  -- 01831: MOV_9
    "11110000",
    "10100100",  -- 01833: MUL
    "00101010",  -- 01834: ADD_1
    "11111010",  -- 01835: MOV_5
    "11101011",  -- 01836: MOV_1
    "00110101",  -- 01837: ADDC_2
    "11110000",
    "11111011",  -- 01839: MOV_5
    "11100100",  -- 01840: CLR_1
    "00111100",  -- 01841: ADDC_1
    "11111100",  -- 01842: MOV_5
    "11101101",  -- 01843: MOV_1
    "10001111",  -- 01844: MOV_9
    "11110000",
    "10100100",  -- 01846: MUL
    "00101011",  -- 01847: ADD_1
    "11111011",  -- 01848: MOV_5
    "11101100",  -- 01849: MOV_1
    "00110101",  -- 01850: ADDC_2
    "11110000",
    "11111100",  -- 01852: MOV_5
    "00100000",  -- 01853: JB
    "11100111",
    "00000011",
    "00010010",  -- 01856: LCALL
    "00000111",
    "10110111",
    "00000010",  -- 01859: LJMP
    "00000101",
    "00110111",
    "10101010",  -- 01862: MOV_6
    "10000010",
    "10101011",  -- 01864: MOV_6
    "10000011",
    "10100010",  -- 01866: MOV_16
    "11110111",
    "00110011",  -- 01868: RLC
    "10010010",  -- 01869: MOV_17
    "11010001",
    "11110101",  -- 01871: MOV_8
    "10000010",
    "01100000",  -- 01873: JZ
    "00000010",
    "11010010",  -- 01875: SETB_2
    "11110111",
    "10101100",  -- 01877: MOV_6
    "11110000",
    "11100101",  -- 01879: MOV_2
    "10000001",
    "00100100",  -- 01881: ADD_4
    "11111001",
    "11111000",  -- 01883: MOV_5
    "11100110",  -- 01884: MOV_3
    "11111101",  -- 01885: MOV_5
    "00001000",  -- 01886: INC_2
    "11100110",  -- 01887: MOV_3
    "11111110",  -- 01888: MOV_5
    "00001000",  -- 01889: INC_2
    "10000110",  -- 01890: MOV_11
    "11110000",
    "00001000",  -- 01892: INC_2
    "11100110",  -- 01893: MOV_3
    "10100010",  -- 01894: MOV_16
    "11110111",
    "00110011",  -- 01896: RLC
    "10010010",  -- 01897: MOV_17
    "11010101",
    "11110101",  -- 01899: MOV_8
    "10000011",
    "01100000",  -- 01901: JZ
    "00000010",
    "11010010",  -- 01903: SETB_2
    "11110111",
    "10101111",  -- 01905: MOV_6
    "11110000",
    "00100010",  -- 01907: RET
    "01100000",  -- 01908: JZ
    "01000000",
    "11111000",  -- 01910: MOV_5
    "00100101",  -- 01911: ADD_2
    "10000010",
    "01010000",  -- 01913: JNC
    "00000010",
    "01110100",  -- 01915: MOV_4
    "11111111",
    "11110101",  -- 01917: MOV_8
    "10000010",
    "11101000",  -- 01919: MOV_1
    "00100100",  -- 01920: ADD_4
    "11111000",
    "01010000",  -- 01922: JNC
    "00011110",
    "11001100",  -- 01924: XCH_1
    "11001011",  -- 01925: XCH_1
    "11001010",  -- 01926: XCH_1
    "11111001",  -- 01927: MOV_5
    "11100100",  -- 01928: CLR_1
    "11001100",  -- 01929: XCH_1
    "00100100",  -- 01930: ADD_4
    "11111000",
    "01010000",  -- 01932: JNC
    "00010100",
    "11001011",  -- 01934: XCH_1
    "11001010",  -- 01935: XCH_1
    "11111001",  -- 01936: MOV_5
    "11100100",  -- 01937: CLR_1
    "11001011",  -- 01938: XCH_1
    "00100100",  -- 01939: ADD_4
    "11111000",
    "01010000",  -- 01941: JNC
    "00001011",
    "11001010",  -- 01943: XCH_1
    "11111001",  -- 01944: MOV_5
    "11100100",  -- 01945: CLR_1
    "11001010",  -- 01946: XCH_1
    "00100100",  -- 01947: ADD_4
    "11111000",
    "01010000",  -- 01949: JNC
    "00000011",
    "01111001",  -- 01951: MOV_7
    "00000000",
    "00100010",  -- 01953: RET
    "00100100",  -- 01954: ADD_4
    "00001000",
    "01100000",  -- 01956: JZ
    "00010000",
    "11111000",  -- 01958: MOV_5
    "11000011",  -- 01959: CLR_2
    "11101100",  -- 01960: MOV_1
    "00010011",  -- 01961: RRC
    "11111100",  -- 01962: MOV_5
    "11101011",  -- 01963: MOV_1
    "00010011",  -- 01964: RRC
    "11111011",  -- 01965: MOV_5
    "11101010",  -- 01966: MOV_1
    "00010011",  -- 01967: RRC
    "11111010",  -- 01968: MOV_5
    "11101001",  -- 01969: MOV_1
    "00010011",  -- 01970: RRC
    "11111001",  -- 01971: MOV_5
    "11011000",  -- 01972: DJNZ_1
    "11110001",
    "00100010",  -- 01974: RET
    "01111000",  -- 01975: MOV_7
    "00000100",
    "11101100",  -- 01977: MOV_1
    "01110000",  -- 01978: JNZ
    "00010001",
    "11100101",  -- 01980: MOV_2
    "10000010",
    "00100100",  -- 01982: ADD_4
    "11111000",
    "01010000",  -- 01984: JNC
    "00001010",
    "11110101",  -- 01986: MOV_8
    "10000010",
    "11100100",  -- 01988: CLR_1
    "11001001",  -- 01989: XCH_1
    "11001010",  -- 01990: XCH_1
    "11001011",  -- 01991: XCH_1
    "11111100",  -- 01992: MOV_5
    "11011000",  -- 01993: DJNZ_1
    "11101111",
    "00100010",  -- 01995: RET
    "11101100",  -- 01996: MOV_1
    "01111000",  -- 01997: MOV_7
    "00100000",
    "00000101",  -- 01999: INC_3
    "10000010",
    "00100000",  -- 02001: JB
    "11100111",
    "00010011",
    "11010101",  -- 02004: DJNZ_2
    "10000010",
    "00000001",
    "00100010",  -- 02007: RET
    "11000011",  -- 02008: CLR_2
    "11101001",  -- 02009: MOV_1
    "00110011",  -- 02010: RLC
    "11111001",  -- 02011: MOV_5
    "11101010",  -- 02012: MOV_1
    "00110011",  -- 02013: RLC
    "11111010",  -- 02014: MOV_5
    "11101011",  -- 02015: MOV_1
    "00110011",  -- 02016: RLC
    "11111011",  -- 02017: MOV_5
    "11101100",  -- 02018: MOV_1
    "00110011",  -- 02019: RLC
    "11111100",  -- 02020: MOV_5
    "11011000",  -- 02021: DJNZ_1
    "11101010",
    "00010101",  -- 02023: DEC_3
    "10000010",
    "00100010",  -- 02025: RET
    "11111111",  -- 02026: MOV_5
    "10101000",  -- 02027: MOV_6
    "10000001",
    "00011000",  -- 02029: DEC_2
    "00011000",  -- 02030: DEC_2
    "00010010",  -- 02031: LCALL
    "00000100",
    "01110111",
    "00010010",  -- 02034: LCALL
    "00000100",
    "01011001",
    "11101001",  -- 02037: MOV_1
    "01100100",  -- 02038: XRL_4
    "00000001",
    "11110101",  -- 02040: MOV_8
    "10000010",
    "00100010",  -- 02042: RET
    "01111111",  -- 02043: MOV_7
    "10011110",
    "00010010",  -- 02045: LCALL
    "00001000",
    "01000001",
    "00110000",  -- 02048: JNB
    "11010001",
    "00000011",
    "00000010",  -- 02051: LJMP
    "00000101",
    "01011000",
    "11000011",  -- 02054: CLR_2
    "11101111",  -- 02055: MOV_1
    "10010101",  -- 02056: SUBB_2
    "10000010",
    "01010000",  -- 02058: JNC
    "00001001",
    "01110100",  -- 02060: MOV_4
    "11111111",
    "11110101",  -- 02062: MOV_8
    "11110000",
    "11110101",  -- 02064: MOV_8
    "10000011",
    "11110101",  -- 02066: MOV_8
    "10000010",
    "00100010",  -- 02068: RET
    "01111001",  -- 02069: MOV_7
    "00000000",
    "00010010",  -- 02071: LCALL
    "00000111",
    "01110100",
    "10001001",  -- 02074: MOV_9
    "10000010",
    "10001010",  -- 02076: MOV_9
    "10000011",
    "10001011",  -- 02078: MOV_9
    "11110000",
    "11101100",  -- 02080: MOV_1
    "00100010",  -- 02081: RET
    "00100000",  -- 02082: JB
    "11110111",
    "00010001",
    "00110000",  -- 02085: JNB
    "11110110",
    "00010011",
    "10001000",  -- 02088: MOV_9
    "10000011",
    "10101000",  -- 02090: MOV_6
    "10000010",
    "00100000",  -- 02092: JB
    "11110101",
    "00001001",
    "11110110",  -- 02095: MOV_13
    "10101000",  -- 02096: MOV_6
    "10000011",
    "01110101",  -- 02098: MOV_12
    "10000011",
    "00000000",
    "00100010",  -- 02101: RET
    "10000000",  -- 02102: SJMP
    "11111110",
    "11110010",  -- 02104: MOVX_3
    "10000000",  -- 02105: SJMP
    "11110101",
    "11110000",  -- 02107: MOVX_4
    "00100010",  -- 02108: RET
    "01110101",  -- 02109: MOV_12
    "10000010",
    "00000000",
    "00100010",  -- 02112: RET
    "10101010",  -- 02113: MOV_6
    "10000010",
    "10101011",  -- 02115: MOV_6
    "10000011",
    "10100010",  -- 02117: MOV_16
    "11110111",
    "00110011",  -- 02119: RLC
    "10010010",  -- 02120: MOV_17
    "11010001",
    "11110101",  -- 02122: MOV_8
    "10000010",
    "01100000",  -- 02124: JZ
    "00000010",
    "11010010",  -- 02126: SETB_2
    "11110111",
    "10101100",  -- 02128: MOV_6
    "11110000",
    "00100010",  -- 02130: RET
    "00000000",  -- 02131: NOP
    "00000000"   -- 02132: NOP
  );
begin
  process (rst, clk)
  begin
    if (rst = '1') then
      data <= CD_8;
    elsif (clk'event and clk = '1') then
      if (rd = '1' and conv_integer(addr) < 2133) then
        data <= PROGRAM(conv_integer(addr));
      else
        data <= CD_8;
      end if;
    end if;
  end process;
end BEHAVIORAL;
